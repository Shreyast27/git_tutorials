sffsdsd
