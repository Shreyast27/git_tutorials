hi sukhitha
