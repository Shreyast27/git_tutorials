ddsfsfsfs
